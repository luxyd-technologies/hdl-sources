
`ifndef __GENERAL_HEADER_DEFS_NONE__
   `define __GENERAL_HEADER_DEFS_NONE__   
   
   `default_nettype none   
 
 
`endif